module vga_Top	(
 
	input 		  clk,
	input [161:0] color,
	input         rst,

	//////////// VGA //////////
	output		          VGA_BLANK_N,
	output reg	  [7:0]  VGA_B,
	output		          VGA_CLK,
	output reg	  [7:0]  VGA_G,
	output		          VGA_HS,
	output reg	  [7:0]  VGA_R,
	output		          VGA_SYNC_N,
	output		          VGA_VS
);

// ----------------------------------------------------
// BITMAP ROM (unchanged)
// ----------------------------------------------------
wire [17:0] SW_db;  // unused but keeping for now

reg [0:0] bitmap_rom [0:3072];

integer i_init;
initial begin
    // Set all to 0 (off) first
    for (i_init = 0; i_init < 3072; i_init = i_init + 1) begin
        bitmap_rom[i_init] = 1'b0;
    end

bitmap_rom[652] = 1'b1;
bitmap_rom[655] = 1'b1;
bitmap_rom[658] = 1'b1;
bitmap_rom[844] = 1'b1;
bitmap_rom[847] = 1'b1;
bitmap_rom[850] = 1'b1;
bitmap_rom[1036] = 1'b1;
bitmap_rom[1039] = 1'b1;
bitmap_rom[1042] = 1'b1;

bitmap_rom[1282] = 1'b1;
bitmap_rom[1285] = 1'b1;
bitmap_rom[1288] = 1'b1;
bitmap_rom[1292] = 1'b1;
bitmap_rom[1295] = 1'b1;
bitmap_rom[1298] = 1'b1;
bitmap_rom[1302] = 1'b1;
bitmap_rom[1305] = 1'b1;
bitmap_rom[1308] = 1'b1;

bitmap_rom[1312] = 1'b1;
bitmap_rom[1315] = 1'b1;
bitmap_rom[1318] = 1'b1;
bitmap_rom[1474] = 1'b1;
bitmap_rom[1477] = 1'b1;
bitmap_rom[1480] = 1'b1;
bitmap_rom[1484] = 1'b1;
bitmap_rom[1487] = 1'b1;
bitmap_rom[1490] = 1'b1;
bitmap_rom[1494] = 1'b1;
bitmap_rom[1497] = 1'b1;
bitmap_rom[1500] = 1'b1;
bitmap_rom[1504] = 1'b1;
bitmap_rom[1507] = 1'b1;
bitmap_rom[1510] = 1'b1;

bitmap_rom[1666] = 1'b1;
bitmap_rom[1669] = 1'b1;
bitmap_rom[1672] = 1'b1;
bitmap_rom[1676] = 1'b1;
bitmap_rom[1679] = 1'b1;
bitmap_rom[1682] = 1'b1;
bitmap_rom[1686] = 1'b1;
bitmap_rom[1689] = 1'b1;
bitmap_rom[1692] = 1'b1;
bitmap_rom[1696] = 1'b1;
bitmap_rom[1699] = 1'b1;
bitmap_rom[1702] = 1'b1;

bitmap_rom[1932] = 1'b1;
bitmap_rom[1935] = 1'b1;
bitmap_rom[1938] = 1'b1;
bitmap_rom[2124] = 1'b1;
bitmap_rom[2127] = 1'b1;
bitmap_rom[2130] = 1'b1;
bitmap_rom[2316] = 1'b1;
bitmap_rom[2319] = 1'b1;
bitmap_rom[2322] = 1'b1;




end

// ----------------------------------------------------
// VGA DRIVER
// ----------------------------------------------------
wire active_pixels;
wire frame_done;
wire [9:0] x;  // current x
wire [9:0] y;  // current y

vga_driver the_vga(
    .clk(clk),
    .rst(rst),

    .vga_clk(VGA_CLK),
    .hsync(VGA_HS),
    .vsync(VGA_VS),

    .active_pixels(active_pixels),
    .frame_done(frame_done),

    .xPixel(x),
    .yPixel(y),

    .VGA_BLANK_N(VGA_BLANK_N),
    .VGA_SYNC_N(VGA_SYNC_N)
);

// ----------------------------------------------------
// MINI FRAMEBUFFER
// ----------------------------------------------------
reg  [14:0] frame_buf_mem_address;
reg  [23:0] frame_buf_mem_data;
reg         frame_buf_mem_wren;
wire [23:0] frame_buf_mem_q;

vga_frame vga_memory(
    .address (frame_buf_mem_address),
    .clock   (clk),
    .data    (frame_buf_mem_data),
    .wren    (frame_buf_mem_wren),
    .q       (frame_buf_mem_q)
);

// ----------------------------------------------------
// FSM + INDEXING
// ----------------------------------------------------
reg [15:0] i;        // loop index for bitmap / framebuffer
reg [7:0]  j;        // bit index into `color` (3 bits per sticker)
reg        blkx;     // indicates whether previous bitmap cell was OFF
reg [7:0]  S, NS;
reg [2:0] write_substate;


parameter 
    START        = 8'd0,
    W2M_INIT     = 8'd1,
    W2M_COND     = 8'd2,
    W2M_INC      = 8'd3,
    RFM_INIT     = 8'd4,
    RFM_DRAWING  = 8'd5,
    ERROR        = 8'hFF;

parameter LOOP_SIZE        = 16'd3072;
parameter LOOP_I_SIZE      = 16'd64;
parameter LOOP_Y_SIZE      = 16'd48;
parameter WIDTH            = 16'd640;
parameter HEIGHT           = 16'd480;
parameter PIXELS_IN_WIDTH  = WIDTH/LOOP_I_SIZE;   // 160
parameter PIXELS_IN_HEIGHT = HEIGHT/LOOP_Y_SIZE;  // 120

// ----------------------------------------------------
// NEXT STATE LOGIC
// ----------------------------------------------------
always @(*) begin
    case (S)
        START:      NS = W2M_INIT;
        W2M_INIT:   NS = W2M_COND;

        W2M_COND: begin
            if (i < LOOP_SIZE)
                NS = W2M_INC;
            else
                NS = RFM_INIT;
        end

        W2M_INC: NS = W2M_COND;

        // After a frame is done, go refresh framebuffer again
        RFM_INIT: begin
            if (frame_done == 1'b1)
                NS = W2M_INIT;
            else
                NS = RFM_INIT;
        end

        RFM_DRAWING: begin
            if (frame_done == 1'b1)
                NS = W2M_INIT;
            else
                NS = RFM_DRAWING;
        end

        default:    NS = ERROR;
    endcase
end

// ----------------------------------------------------
// STATE REGISTER
// ----------------------------------------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        S  <= START;
    end else begin
        S  <= NS;
    end
end

// ----------------------------------------------------
// SEQUENTIAL: WRITE/READ CONTROL + j / blkx UPDATE
// ----------------------------------------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        frame_buf_mem_address <= 14'd0;
        frame_buf_mem_data    <= 24'd0;
        frame_buf_mem_wren    <= 1'b0;
        i                     <= 16'd0;
        j                     <= 8'd0;
		  write_substate <= 3'b000;
    end else begin
        case (S)
            START: begin
                frame_buf_mem_address <= 14'd0;
                frame_buf_mem_data    <= 24'd0;
                frame_buf_mem_wren    <= 1'b0;
                i                     <= 16'd0;
                j                     <= 8'd0;
					 write_substate <= 3'b000;
            end

            // Start a new write pass
            W2M_INIT: begin
                frame_buf_mem_address <= 14'd0;
                frame_buf_mem_data    <= 24'd0;
                frame_buf_mem_wren    <= 1'b1;
                i                     <= 16'd0;
                j                     <= 8'd0;  
					write_substate <= 3'b000; // restart color bit index
            end

            W2M_COND: begin
                // nothing to do here; controlled by NS logic
            end

            // Write one pixel's worth of RGB to the framebuffer
            W2M_INC: begin
    if (bitmap_rom[i] == 1'b1) begin
        case (write_substate)
            3'b000: begin
                frame_buf_mem_address <= i;
                frame_buf_mem_data    <= {red, green, blue};
                write_substate        <= 3'b001;
            end

            3'b001: begin
                frame_buf_mem_address <= i + 1;
                frame_buf_mem_data    <= {red, green, blue};
                write_substate        <= 3'b010;
            end

            3'b010: begin
                frame_buf_mem_address <= i + LOOP_I_SIZE;  // = +64
                frame_buf_mem_data    <= {red, green, blue};
                write_substate        <= 3'b011;
            end

            3'b011: begin
                frame_buf_mem_address <= i + LOOP_I_SIZE + 1; // = +65
                frame_buf_mem_data    <= {red, green, blue};
                write_substate        <= 3'b100;
            end

            3'b100: begin
                // done writing this 2×2 block
                i <= i + 1;
                j <= j + 3;
                write_substate <= 3'b000;
            end
        endcase
    end else begin
        // OFF pixel: skip writing
        i <= i + 1;
    end
end
            // Read phase: map x/y to framebuffer address
            RFM_INIT: begin
                frame_buf_mem_wren <= 1'b0; // turn off writing
                if (y < HEIGHT && x < WIDTH)
                    frame_buf_mem_address <= (y/PIXELS_IN_HEIGHT) * LOOP_I_SIZE + (x/PIXELS_IN_WIDTH);
            end

            RFM_DRAWING: begin
                if (y < HEIGHT && x < WIDTH)
                    frame_buf_mem_address <= (y/PIXELS_IN_HEIGHT) * LOOP_I_SIZE + (x/PIXELS_IN_WIDTH);
            end

            default: begin
                // do nothing
            end
        endcase
    end
end

// ----------------------------------------------------
// COMBINATIONAL: COLOR MAPPING (NO STATE UPDATES)
// ----------------------------------------------------
reg [7:0] red;
reg [7:0] green;
reg [7:0] blue;
reg [2:0] packedColor;

always @(*) begin
    // Always show what's in memory on the VGA outputs
    {VGA_R, VGA_G, VGA_B} = frame_buf_mem_q;

    // Default RGB if bitmap cell is OFF
    red   = 8'h00;
    green = 8'h00;
    blue  = 8'h00;
    packedColor = 3'b000;

    // Only compute a color when we're in the write phase and the bitmap cell is ON
    // (During read phase, `red/green/blue` only matter indirectly via previous W2M pass).
    if (bitmap_rom[i] == 1'b1) begin
        // NOTE: j points to the *current* sticker's 3-bit color in `color`.
        packedColor[0] = color[j];
        packedColor[1] = color[j+1];
        packedColor[2] = color[j+2];

        // Map 3-bit packedColor to RGB
        if      (packedColor == 3'b000) begin
            red   = 8'hFF;
            green = 8'hFF;
            blue  = 8'hFF;
        end else if (packedColor == 3'b001) begin
            red   = 8'hFF;
            green = 8'h40;
            blue  = 8'h00;
        end else if (packedColor == 3'b010) begin
            red   = 8'h00;
            green = 8'hFF;
            blue  = 8'h00;
        end else if (packedColor == 3'b011) begin
            red   = 8'hFF;
            green = 8'h00;
            blue  = 8'h00;
        end else if (packedColor == 3'b100) begin
            red   = 8'h00;
            green = 8'h00;
            blue  = 8'hFF;
        end else if (packedColor == 3'b101) begin
            red   = 8'hFF;
            green = 8'hFF;
            blue  = 8'h00;
        end else begin
            // fallback / error color (magenta)
            red   = 8'hFF;
            green = 8'h00;
            blue  = 8'hFF;
        end
    end
end

endmodule